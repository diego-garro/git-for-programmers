module main

fn main() {
	println('Hello World!')
	println('I just added this in VSCode')
	println('This line added to show the staging area')
}
