module main

import time

fn main() {
	println('Hello World!')
	println('I just added this in VSCode')
	println('This line added to show the staging area')
}

struct Book {
	pub:
		title string
		authors string[]
		publication_date time.Time
}
