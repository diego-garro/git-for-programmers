module main

fn main() {
	println('Hello World!')
	println('I just added this in VSCode')
}
